module top_module( input in, output out );

	assign out = in; // continuous assignment --> the value of in will be driven to out whenever a value is drivien to in
    
endmodule